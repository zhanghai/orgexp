`timescale 1ns / 1ps

module Decode_pc_Int(
		input clk,
		input reset,
		input INT,
		input RFE,
		input [31:0] pc_next,
		output reg [31:0] pc
		);
endmodule
