`timescale 1ns / 1ps

module clk_div(
		input clk,
		input rst,
		input SW2,
		output [31:0] clkdiv,
		output Clk_CPU
		);
endmodule
